****comparator test*****

X1 1 1d 0 v_p v_n Vout comparatorP

*****************************************
.include osu018.lib
******************************************


***********ComparatorLOW******************


.subckt comparatorP N001 N002 0 vp vn Vout
ME1 N003 N004 N001 N001 pfet l=200n w=2u m=1
*ME2 N004 N004 N001 N001 pfet l=200n w=2u m=1
ME2 N004 N004 0 0 nfet l=200n w=2u m=1

M1 N005 vn N003 N001 pfet l=200n w=2u m=1
M2 N006 vp N003 N001 pfet l=200n w=2u m=1
M3 N005 N005 0 0 nfet l=200n w=2u m=1
M4 N006 N005 0 0 nfet l=200n w=2u m=1
M5 N007 N004 N001 N001 pfet l=200n w=2u m=1
M6 N007 N006 0 0 nfet l=200n w=6u m=1
M8 N008 N007 N002 N002 pfet l=200n w=1u
M9 Vout N008 N002 N002 pfet l=200n w=1u
M10 N008 N007 0 0 nfet l=200n w=5u
M11 Vout N008 0 0 nfet l=200n w=5u
R N001 N004 50k
.ends comparatorP


************************************

*************************************

V_a 1 0 pulse(0 3.3 1n 1n 1n 3u 6u)
V_d 1d 0 3.3V


Vp v_p 0 pulse(0.408v 0.4v 1n 1n 1n 1u 2u)
Vn v_n 0 pulse(0.4v 0.408v 1n 1n 1n 1u 2u)



*************************************
.tran 1ns 6us
.control

run
plot V(v_p)+0.01 V(v_n)
plot V(Vout)+4 V(1)
.endc
.end




