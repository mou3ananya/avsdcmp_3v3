magic
tech scmos
timestamp 1599951872
<< nwell >>
rect -210 78 -64 158
rect -58 105 26 146
rect 32 117 132 158
rect -58 63 -4 105
rect 84 101 132 117
rect -67 -56 12 24
rect 26 23 78 63
<< ntransistor >>
rect -196 45 -194 65
rect -175 45 -173 65
rect -122 50 -120 60
rect -101 50 -99 60
rect -80 50 -78 60
rect -41 37 -39 57
rect -20 37 -18 57
rect 10 37 12 97
rect 47 89 49 99
rect 68 89 70 99
rect 99 59 101 69
rect 107 59 109 69
rect 115 59 117 69
rect -212 -108 -210 -8
rect -180 -22 -178 -2
rect -159 -22 -157 -2
rect 41 -5 43 5
rect 62 -5 64 5
rect -53 -89 -51 -69
rect -32 -89 -30 -69
rect -37 -146 -35 -126
rect -16 -146 -14 -126
<< ptransistor >>
rect -196 87 -194 107
rect -175 87 -173 107
rect -147 87 -145 147
rect -122 85 -120 105
rect -101 85 -99 105
rect -80 85 -78 105
rect -32 102 -30 122
rect 10 111 12 131
rect 47 124 49 144
rect 68 124 70 144
rect 99 107 101 147
rect 104 107 106 147
rect 112 127 114 147
rect -41 69 -39 89
rect -20 69 -18 89
rect 41 30 43 50
rect 62 30 64 50
rect -53 -47 -51 -27
rect -32 -47 -30 -27
rect -4 -47 -2 13
<< ndiffusion >>
rect 2 93 3 97
rect 7 93 10 97
rect 2 92 10 93
rect -204 61 -203 65
rect -199 61 -196 65
rect -204 60 -196 61
rect -204 56 -203 60
rect -199 56 -196 60
rect -204 55 -196 56
rect -204 51 -203 55
rect -199 51 -196 55
rect -204 50 -196 51
rect -204 46 -203 50
rect -199 46 -196 50
rect -204 45 -196 46
rect -194 64 -186 65
rect -194 60 -191 64
rect -187 60 -186 64
rect -194 59 -186 60
rect -194 55 -191 59
rect -187 55 -186 59
rect -194 54 -186 55
rect -194 50 -191 54
rect -187 50 -186 54
rect -194 49 -186 50
rect -194 45 -191 49
rect -187 45 -186 49
rect -183 61 -182 65
rect -178 61 -175 65
rect -183 60 -175 61
rect -183 56 -182 60
rect -178 56 -175 60
rect -183 55 -175 56
rect -183 51 -182 55
rect -178 51 -175 55
rect -183 50 -175 51
rect -183 46 -182 50
rect -178 46 -175 50
rect -183 45 -175 46
rect -173 64 -165 65
rect -173 60 -170 64
rect -166 60 -165 64
rect 2 88 3 92
rect 7 88 10 92
rect 2 87 10 88
rect 2 83 3 87
rect 7 83 10 87
rect 2 82 10 83
rect 2 78 3 82
rect 7 78 10 82
rect 2 77 10 78
rect 2 73 3 77
rect 7 73 10 77
rect 2 72 10 73
rect 2 68 3 72
rect 7 68 10 72
rect 2 67 10 68
rect 2 63 3 67
rect 7 63 10 67
rect 2 62 10 63
rect -173 59 -165 60
rect -173 55 -170 59
rect -166 55 -165 59
rect -173 54 -165 55
rect -173 50 -170 54
rect -166 50 -165 54
rect -130 56 -129 60
rect -125 56 -122 60
rect -130 55 -122 56
rect -130 51 -129 55
rect -125 51 -122 55
rect -130 50 -122 51
rect -120 59 -112 60
rect -120 55 -117 59
rect -113 55 -112 59
rect -120 54 -112 55
rect -120 50 -117 54
rect -113 50 -112 54
rect -109 56 -108 60
rect -104 56 -101 60
rect -109 55 -101 56
rect -109 51 -108 55
rect -104 51 -101 55
rect -109 50 -101 51
rect -99 59 -91 60
rect -99 55 -96 59
rect -92 55 -91 59
rect -99 54 -91 55
rect -99 50 -96 54
rect -92 50 -91 54
rect -88 56 -87 60
rect -83 56 -80 60
rect -88 55 -80 56
rect -88 51 -87 55
rect -83 51 -80 55
rect -88 50 -80 51
rect -78 59 -70 60
rect -78 55 -75 59
rect -71 55 -70 59
rect 2 58 3 62
rect 7 58 10 62
rect 2 57 10 58
rect -78 54 -70 55
rect -78 50 -75 54
rect -71 50 -70 54
rect -49 53 -48 57
rect -44 53 -41 57
rect -49 52 -41 53
rect -173 49 -165 50
rect -173 45 -170 49
rect -166 45 -165 49
rect -49 48 -48 52
rect -44 48 -41 52
rect -49 47 -41 48
rect -49 43 -48 47
rect -44 43 -41 47
rect -49 42 -41 43
rect -49 38 -48 42
rect -44 38 -41 42
rect -49 37 -41 38
rect -39 56 -31 57
rect -39 52 -36 56
rect -32 52 -31 56
rect -39 51 -31 52
rect -39 47 -36 51
rect -32 47 -31 51
rect -39 46 -31 47
rect -39 42 -36 46
rect -32 42 -31 46
rect -39 41 -31 42
rect -39 37 -36 41
rect -32 37 -31 41
rect -28 55 -20 57
rect -28 51 -27 55
rect -23 51 -20 55
rect -28 50 -20 51
rect -28 46 -27 50
rect -23 46 -20 50
rect -28 45 -20 46
rect -28 41 -27 45
rect -23 41 -20 45
rect -28 37 -20 41
rect -18 56 -10 57
rect -18 52 -15 56
rect -11 52 -10 56
rect -18 51 -10 52
rect -18 47 -15 51
rect -11 47 -10 51
rect -18 46 -10 47
rect -18 42 -15 46
rect -11 42 -10 46
rect -18 41 -10 42
rect -18 37 -15 41
rect -11 37 -10 41
rect 2 53 3 57
rect 7 53 10 57
rect 2 52 10 53
rect 2 48 3 52
rect 7 48 10 52
rect 2 47 10 48
rect 2 43 3 47
rect 7 43 10 47
rect 2 42 10 43
rect 2 38 3 42
rect 7 38 10 42
rect 2 37 10 38
rect 12 96 20 97
rect 12 92 15 96
rect 19 92 20 96
rect 12 91 20 92
rect 12 87 15 91
rect 19 87 20 91
rect 39 95 40 99
rect 44 95 47 99
rect 39 94 47 95
rect 39 90 40 94
rect 44 90 47 94
rect 39 89 47 90
rect 49 98 57 99
rect 49 94 52 98
rect 56 94 57 98
rect 49 93 57 94
rect 49 89 52 93
rect 56 89 57 93
rect 60 95 61 99
rect 65 95 68 99
rect 60 94 68 95
rect 60 90 61 94
rect 65 90 68 94
rect 60 89 68 90
rect 70 98 78 99
rect 70 94 73 98
rect 77 94 78 98
rect 70 93 78 94
rect 70 89 73 93
rect 77 89 78 93
rect 12 86 20 87
rect 12 82 15 86
rect 19 82 20 86
rect 12 81 20 82
rect 12 77 15 81
rect 19 77 20 81
rect 12 76 20 77
rect 12 72 15 76
rect 19 72 20 76
rect 12 71 20 72
rect 12 67 15 71
rect 19 67 20 71
rect 12 66 20 67
rect 12 62 15 66
rect 19 62 20 66
rect 12 61 20 62
rect 12 57 15 61
rect 19 57 20 61
rect 12 56 20 57
rect 98 59 99 69
rect 101 59 102 69
rect 106 59 107 69
rect 109 59 110 69
rect 114 59 115 69
rect 117 59 118 69
rect 12 52 15 56
rect 19 52 20 56
rect 12 51 20 52
rect 12 47 15 51
rect 19 47 20 51
rect 12 46 20 47
rect 12 42 15 46
rect 19 42 20 46
rect 12 41 20 42
rect 12 37 15 41
rect 19 37 20 41
rect -188 -6 -187 -2
rect -183 -6 -180 -2
rect -188 -7 -180 -6
rect -220 -12 -219 -8
rect -215 -12 -212 -8
rect -220 -13 -212 -12
rect -220 -17 -219 -13
rect -215 -17 -212 -13
rect -220 -18 -212 -17
rect -220 -22 -219 -18
rect -215 -22 -212 -18
rect -220 -23 -212 -22
rect -220 -27 -219 -23
rect -215 -27 -212 -23
rect -220 -28 -212 -27
rect -220 -32 -219 -28
rect -215 -32 -212 -28
rect -220 -33 -212 -32
rect -220 -37 -219 -33
rect -215 -37 -212 -33
rect -220 -38 -212 -37
rect -220 -42 -219 -38
rect -215 -42 -212 -38
rect -220 -43 -212 -42
rect -220 -47 -219 -43
rect -215 -47 -212 -43
rect -220 -48 -212 -47
rect -220 -52 -219 -48
rect -215 -52 -212 -48
rect -220 -53 -212 -52
rect -220 -57 -219 -53
rect -215 -57 -212 -53
rect -220 -58 -212 -57
rect -220 -62 -219 -58
rect -215 -62 -212 -58
rect -220 -63 -212 -62
rect -220 -67 -219 -63
rect -215 -67 -212 -63
rect -220 -68 -212 -67
rect -220 -72 -219 -68
rect -215 -72 -212 -68
rect -220 -73 -212 -72
rect -220 -77 -219 -73
rect -215 -77 -212 -73
rect -220 -78 -212 -77
rect -220 -82 -219 -78
rect -215 -82 -212 -78
rect -220 -83 -212 -82
rect -220 -87 -219 -83
rect -215 -87 -212 -83
rect -220 -88 -212 -87
rect -220 -92 -219 -88
rect -215 -92 -212 -88
rect -220 -93 -212 -92
rect -220 -97 -219 -93
rect -215 -97 -212 -93
rect -220 -98 -212 -97
rect -220 -102 -219 -98
rect -215 -102 -212 -98
rect -220 -103 -212 -102
rect -220 -107 -219 -103
rect -215 -107 -212 -103
rect -220 -108 -212 -107
rect -210 -9 -202 -8
rect -210 -13 -207 -9
rect -203 -13 -202 -9
rect -210 -14 -202 -13
rect -210 -18 -207 -14
rect -203 -18 -202 -14
rect -210 -19 -202 -18
rect -210 -23 -207 -19
rect -203 -23 -202 -19
rect -188 -11 -187 -7
rect -183 -11 -180 -7
rect -188 -12 -180 -11
rect -188 -16 -187 -12
rect -183 -16 -180 -12
rect -188 -17 -180 -16
rect -188 -21 -187 -17
rect -183 -21 -180 -17
rect -188 -22 -180 -21
rect -178 -3 -170 -2
rect -178 -7 -175 -3
rect -171 -7 -170 -3
rect -178 -8 -170 -7
rect -178 -12 -175 -8
rect -171 -12 -170 -8
rect -178 -13 -170 -12
rect -178 -17 -175 -13
rect -171 -17 -170 -13
rect -178 -18 -170 -17
rect -178 -22 -175 -18
rect -171 -22 -170 -18
rect -167 -6 -166 -2
rect -162 -6 -159 -2
rect -167 -7 -159 -6
rect -167 -11 -166 -7
rect -162 -11 -159 -7
rect -167 -12 -159 -11
rect -167 -16 -166 -12
rect -162 -16 -159 -12
rect -167 -17 -159 -16
rect -167 -21 -166 -17
rect -162 -21 -159 -17
rect -167 -22 -159 -21
rect -157 -3 -149 -2
rect -157 -7 -154 -3
rect -150 -7 -149 -3
rect -157 -8 -149 -7
rect -157 -12 -154 -8
rect -150 -12 -149 -8
rect -157 -13 -149 -12
rect -157 -17 -154 -13
rect -150 -17 -149 -13
rect -157 -18 -149 -17
rect -157 -22 -154 -18
rect -150 -22 -149 -18
rect -210 -24 -202 -23
rect -210 -28 -207 -24
rect -203 -28 -202 -24
rect -210 -29 -202 -28
rect -210 -33 -207 -29
rect -203 -33 -202 -29
rect -210 -34 -202 -33
rect -210 -38 -207 -34
rect -203 -38 -202 -34
rect -210 -39 -202 -38
rect -210 -43 -207 -39
rect -203 -43 -202 -39
rect -210 -44 -202 -43
rect -210 -48 -207 -44
rect -203 -48 -202 -44
rect 33 1 34 5
rect 38 1 41 5
rect 33 0 41 1
rect 33 -4 34 0
rect 38 -4 41 0
rect 33 -5 41 -4
rect 43 4 51 5
rect 43 0 46 4
rect 50 0 51 4
rect 43 -1 51 0
rect 43 -5 46 -1
rect 50 -5 51 -1
rect 54 1 55 5
rect 59 1 62 5
rect 54 0 62 1
rect 54 -4 55 0
rect 59 -4 62 0
rect 54 -5 62 -4
rect 64 4 72 5
rect 64 0 67 4
rect 71 0 72 4
rect 64 -1 72 0
rect 64 -5 67 -1
rect 71 -5 72 -1
rect -210 -49 -202 -48
rect -210 -53 -207 -49
rect -203 -53 -202 -49
rect -210 -54 -202 -53
rect -210 -58 -207 -54
rect -203 -58 -202 -54
rect -210 -59 -202 -58
rect -210 -63 -207 -59
rect -203 -63 -202 -59
rect -210 -64 -202 -63
rect -210 -68 -207 -64
rect -203 -68 -202 -64
rect -210 -69 -202 -68
rect -210 -73 -207 -69
rect -203 -73 -202 -69
rect -210 -74 -202 -73
rect -210 -78 -207 -74
rect -203 -78 -202 -74
rect -210 -79 -202 -78
rect -210 -83 -207 -79
rect -203 -83 -202 -79
rect -210 -84 -202 -83
rect -210 -88 -207 -84
rect -203 -88 -202 -84
rect -210 -89 -202 -88
rect -61 -73 -60 -69
rect -56 -73 -53 -69
rect -61 -74 -53 -73
rect -61 -78 -60 -74
rect -56 -78 -53 -74
rect -61 -79 -53 -78
rect -61 -83 -60 -79
rect -56 -83 -53 -79
rect -61 -84 -53 -83
rect -61 -88 -60 -84
rect -56 -88 -53 -84
rect -61 -89 -53 -88
rect -51 -70 -43 -69
rect -51 -74 -48 -70
rect -44 -74 -43 -70
rect -51 -75 -43 -74
rect -51 -79 -48 -75
rect -44 -79 -43 -75
rect -51 -80 -43 -79
rect -51 -84 -48 -80
rect -44 -84 -43 -80
rect -51 -85 -43 -84
rect -51 -89 -48 -85
rect -44 -89 -43 -85
rect -40 -73 -39 -69
rect -35 -73 -32 -69
rect -40 -74 -32 -73
rect -40 -78 -39 -74
rect -35 -78 -32 -74
rect -40 -79 -32 -78
rect -40 -83 -39 -79
rect -35 -83 -32 -79
rect -40 -84 -32 -83
rect -40 -88 -39 -84
rect -35 -88 -32 -84
rect -40 -89 -32 -88
rect -30 -70 -22 -69
rect -30 -74 -27 -70
rect -23 -74 -22 -70
rect -30 -75 -22 -74
rect -30 -79 -27 -75
rect -23 -79 -22 -75
rect -30 -80 -22 -79
rect -30 -84 -27 -80
rect -23 -84 -22 -80
rect -30 -85 -22 -84
rect -30 -89 -27 -85
rect -23 -89 -22 -85
rect -210 -93 -207 -89
rect -203 -93 -202 -89
rect -210 -94 -202 -93
rect -210 -98 -207 -94
rect -203 -98 -202 -94
rect -210 -99 -202 -98
rect -210 -103 -207 -99
rect -203 -103 -202 -99
rect -210 -104 -202 -103
rect -210 -108 -207 -104
rect -203 -108 -202 -104
rect -45 -130 -44 -126
rect -40 -130 -37 -126
rect -45 -131 -37 -130
rect -45 -135 -44 -131
rect -40 -135 -37 -131
rect -45 -136 -37 -135
rect -45 -140 -44 -136
rect -40 -140 -37 -136
rect -45 -141 -37 -140
rect -45 -145 -44 -141
rect -40 -145 -37 -141
rect -45 -146 -37 -145
rect -35 -127 -27 -126
rect -35 -131 -32 -127
rect -28 -131 -27 -127
rect -35 -132 -27 -131
rect -35 -136 -32 -132
rect -28 -136 -27 -132
rect -35 -137 -27 -136
rect -35 -141 -32 -137
rect -28 -141 -27 -137
rect -35 -142 -27 -141
rect -35 -146 -32 -142
rect -28 -146 -27 -142
rect -24 -130 -23 -126
rect -19 -130 -16 -126
rect -24 -131 -16 -130
rect -24 -135 -23 -131
rect -19 -135 -16 -131
rect -24 -136 -16 -135
rect -24 -140 -23 -136
rect -19 -140 -16 -136
rect -24 -141 -16 -140
rect -24 -145 -23 -141
rect -19 -145 -16 -141
rect -24 -146 -16 -145
rect -14 -127 -6 -126
rect -14 -131 -11 -127
rect -7 -131 -6 -127
rect -14 -132 -6 -131
rect -14 -136 -11 -132
rect -7 -136 -6 -132
rect -14 -137 -6 -136
rect -14 -141 -11 -137
rect -7 -141 -6 -137
rect -14 -142 -6 -141
rect -14 -146 -11 -142
rect -7 -146 -6 -142
<< pdiffusion >>
rect -155 146 -147 147
rect -155 142 -154 146
rect -150 142 -147 146
rect -155 141 -147 142
rect -155 137 -154 141
rect -150 137 -147 141
rect -155 136 -147 137
rect -155 132 -154 136
rect -150 132 -147 136
rect -155 131 -147 132
rect -155 127 -154 131
rect -150 127 -147 131
rect -155 126 -147 127
rect -155 122 -154 126
rect -150 122 -147 126
rect -155 121 -147 122
rect -155 117 -154 121
rect -150 117 -147 121
rect -155 116 -147 117
rect -155 112 -154 116
rect -150 112 -147 116
rect -155 111 -147 112
rect -155 107 -154 111
rect -150 107 -147 111
rect -204 106 -196 107
rect -204 102 -203 106
rect -199 102 -196 106
rect -204 101 -196 102
rect -204 97 -203 101
rect -199 97 -196 101
rect -204 96 -196 97
rect -204 92 -203 96
rect -199 92 -196 96
rect -204 91 -196 92
rect -204 87 -203 91
rect -199 87 -196 91
rect -194 103 -191 107
rect -187 103 -186 107
rect -194 102 -186 103
rect -194 98 -191 102
rect -187 98 -186 102
rect -194 97 -186 98
rect -194 93 -191 97
rect -187 93 -186 97
rect -194 92 -186 93
rect -194 88 -191 92
rect -187 88 -186 92
rect -194 87 -186 88
rect -183 106 -175 107
rect -183 102 -182 106
rect -178 102 -175 106
rect -183 101 -175 102
rect -183 97 -182 101
rect -178 97 -175 101
rect -183 96 -175 97
rect -183 92 -182 96
rect -178 92 -175 96
rect -183 91 -175 92
rect -183 87 -182 91
rect -178 87 -175 91
rect -173 103 -170 107
rect -166 103 -165 107
rect -173 102 -165 103
rect -173 98 -170 102
rect -166 98 -165 102
rect -173 97 -165 98
rect -173 93 -170 97
rect -166 93 -165 97
rect -173 92 -165 93
rect -173 88 -170 92
rect -166 88 -165 92
rect -173 87 -165 88
rect -155 106 -147 107
rect -155 102 -154 106
rect -150 102 -147 106
rect -155 101 -147 102
rect -155 97 -154 101
rect -150 97 -147 101
rect -155 96 -147 97
rect -155 92 -154 96
rect -150 92 -147 96
rect -155 91 -147 92
rect -155 87 -154 91
rect -150 87 -147 91
rect -145 143 -142 147
rect -138 143 -137 147
rect 39 143 47 144
rect -145 142 -137 143
rect -145 138 -142 142
rect -138 138 -137 142
rect 39 139 40 143
rect 44 139 47 143
rect -145 137 -137 138
rect -145 133 -142 137
rect -138 133 -137 137
rect 39 138 47 139
rect -145 132 -137 133
rect -145 128 -142 132
rect -138 128 -137 132
rect -145 127 -137 128
rect -145 123 -142 127
rect -138 123 -137 127
rect -145 122 -137 123
rect 39 134 40 138
rect 44 134 47 138
rect 39 133 47 134
rect 2 130 10 131
rect 2 126 3 130
rect 7 126 10 130
rect 2 125 10 126
rect -145 118 -142 122
rect -138 118 -137 122
rect -145 117 -137 118
rect -145 113 -142 117
rect -138 113 -137 117
rect -145 112 -137 113
rect -145 108 -142 112
rect -138 108 -137 112
rect -40 121 -32 122
rect -40 117 -39 121
rect -35 117 -32 121
rect -40 116 -32 117
rect -40 112 -39 116
rect -35 112 -32 116
rect -40 111 -32 112
rect -145 107 -137 108
rect -145 103 -142 107
rect -138 103 -137 107
rect -40 107 -39 111
rect -35 107 -32 111
rect -40 106 -32 107
rect -145 102 -137 103
rect -145 98 -142 102
rect -138 98 -137 102
rect -145 97 -137 98
rect -145 93 -142 97
rect -138 93 -137 97
rect -145 92 -137 93
rect -145 88 -142 92
rect -138 88 -137 92
rect -145 87 -137 88
rect -130 104 -122 105
rect -130 100 -129 104
rect -125 100 -122 104
rect -130 99 -122 100
rect -130 95 -129 99
rect -125 95 -122 99
rect -130 94 -122 95
rect -130 90 -129 94
rect -125 90 -122 94
rect -130 89 -122 90
rect -130 85 -129 89
rect -125 85 -122 89
rect -120 101 -117 105
rect -113 101 -112 105
rect -120 100 -112 101
rect -120 96 -117 100
rect -113 96 -112 100
rect -120 95 -112 96
rect -120 91 -117 95
rect -113 91 -112 95
rect -120 90 -112 91
rect -120 86 -117 90
rect -113 86 -112 90
rect -120 85 -112 86
rect -109 104 -101 105
rect -109 100 -108 104
rect -104 100 -101 104
rect -109 99 -101 100
rect -109 95 -108 99
rect -104 95 -101 99
rect -109 94 -101 95
rect -109 90 -108 94
rect -104 90 -101 94
rect -109 89 -101 90
rect -109 85 -108 89
rect -104 85 -101 89
rect -99 101 -96 105
rect -92 101 -91 105
rect -99 100 -91 101
rect -99 96 -96 100
rect -92 96 -91 100
rect -99 95 -91 96
rect -99 91 -96 95
rect -92 91 -91 95
rect -99 90 -91 91
rect -99 86 -96 90
rect -92 86 -91 90
rect -99 85 -91 86
rect -88 104 -80 105
rect -88 100 -87 104
rect -83 100 -80 104
rect -88 99 -80 100
rect -88 95 -87 99
rect -83 95 -80 99
rect -88 94 -80 95
rect -88 90 -87 94
rect -83 90 -80 94
rect -88 89 -80 90
rect -88 85 -87 89
rect -83 85 -80 89
rect -78 101 -75 105
rect -71 101 -70 105
rect -40 102 -39 106
rect -35 102 -32 106
rect -30 118 -27 122
rect -23 118 -22 122
rect -30 117 -22 118
rect -30 113 -27 117
rect -23 113 -22 117
rect -30 112 -22 113
rect 2 121 3 125
rect 7 121 10 125
rect 2 120 10 121
rect 2 116 3 120
rect 7 116 10 120
rect 2 115 10 116
rect -30 108 -27 112
rect -23 108 -22 112
rect -30 107 -22 108
rect -30 103 -27 107
rect -23 103 -22 107
rect -30 102 -22 103
rect 2 111 3 115
rect 7 111 10 115
rect 12 127 15 131
rect 19 127 20 131
rect 12 126 20 127
rect 12 122 15 126
rect 19 122 20 126
rect 39 129 40 133
rect 44 129 47 133
rect 39 128 47 129
rect 39 124 40 128
rect 44 124 47 128
rect 49 140 52 144
rect 56 140 57 144
rect 49 139 57 140
rect 49 135 52 139
rect 56 135 57 139
rect 49 134 57 135
rect 49 130 52 134
rect 56 130 57 134
rect 49 129 57 130
rect 49 125 52 129
rect 56 125 57 129
rect 49 124 57 125
rect 60 143 68 144
rect 60 139 61 143
rect 65 139 68 143
rect 60 138 68 139
rect 60 134 61 138
rect 65 134 68 138
rect 60 133 68 134
rect 60 129 61 133
rect 65 129 68 133
rect 60 128 68 129
rect 60 124 61 128
rect 65 124 68 128
rect 70 140 73 144
rect 77 140 78 144
rect 70 139 78 140
rect 70 135 73 139
rect 77 135 78 139
rect 70 134 78 135
rect 70 130 73 134
rect 77 130 78 134
rect 70 129 78 130
rect 70 125 73 129
rect 77 125 78 129
rect 70 124 78 125
rect 12 121 20 122
rect 12 117 15 121
rect 19 117 20 121
rect 12 116 20 117
rect 12 112 15 116
rect 19 112 20 116
rect 12 111 20 112
rect -78 100 -70 101
rect -78 96 -75 100
rect -71 96 -70 100
rect -78 95 -70 96
rect -78 91 -75 95
rect -71 91 -70 95
rect -78 90 -70 91
rect -78 86 -75 90
rect -71 86 -70 90
rect 98 107 99 147
rect 101 107 104 147
rect 106 107 107 147
rect 111 127 112 147
rect 114 127 115 147
rect -78 85 -70 86
rect -49 88 -41 89
rect -49 84 -48 88
rect -44 84 -41 88
rect -49 83 -41 84
rect -49 79 -48 83
rect -44 79 -41 83
rect -49 78 -41 79
rect -49 74 -48 78
rect -44 74 -41 78
rect -49 73 -41 74
rect -49 69 -48 73
rect -44 69 -41 73
rect -39 85 -36 89
rect -32 85 -31 89
rect -39 84 -31 85
rect -39 80 -36 84
rect -32 80 -31 84
rect -39 79 -31 80
rect -39 75 -36 79
rect -32 75 -31 79
rect -39 74 -31 75
rect -39 70 -36 74
rect -32 70 -31 74
rect -39 69 -31 70
rect -28 88 -20 89
rect -28 84 -27 88
rect -23 84 -20 88
rect -28 83 -20 84
rect -28 79 -27 83
rect -23 79 -20 83
rect -28 78 -20 79
rect -28 74 -27 78
rect -23 74 -20 78
rect -28 73 -20 74
rect -28 69 -27 73
rect -23 69 -20 73
rect -18 85 -15 89
rect -11 85 -10 89
rect -18 84 -10 85
rect -18 80 -15 84
rect -11 80 -10 84
rect -18 79 -10 80
rect -18 75 -15 79
rect -11 75 -10 79
rect -18 74 -10 75
rect -18 70 -15 74
rect -11 70 -10 74
rect -18 69 -10 70
rect 33 49 41 50
rect 33 45 34 49
rect 38 45 41 49
rect 33 44 41 45
rect 33 40 34 44
rect 38 40 41 44
rect 33 39 41 40
rect 33 35 34 39
rect 38 35 41 39
rect 33 34 41 35
rect 33 30 34 34
rect 38 30 41 34
rect 43 46 46 50
rect 50 46 51 50
rect 43 45 51 46
rect 43 41 46 45
rect 50 41 51 45
rect 43 40 51 41
rect 43 36 46 40
rect 50 36 51 40
rect 43 35 51 36
rect 43 31 46 35
rect 50 31 51 35
rect 43 30 51 31
rect 54 49 62 50
rect 54 45 55 49
rect 59 45 62 49
rect 54 44 62 45
rect 54 40 55 44
rect 59 40 62 44
rect 54 39 62 40
rect 54 35 55 39
rect 59 35 62 39
rect 54 34 62 35
rect 54 30 55 34
rect 59 30 62 34
rect 64 46 67 50
rect 71 46 72 50
rect 64 45 72 46
rect 64 41 67 45
rect 71 41 72 45
rect 64 40 72 41
rect 64 36 67 40
rect 71 36 72 40
rect 64 35 72 36
rect 64 31 67 35
rect 71 31 72 35
rect 64 30 72 31
rect -12 12 -4 13
rect -12 8 -11 12
rect -7 8 -4 12
rect -12 7 -4 8
rect -12 3 -11 7
rect -7 3 -4 7
rect -12 2 -4 3
rect -12 -2 -11 2
rect -7 -2 -4 2
rect -12 -3 -4 -2
rect -12 -7 -11 -3
rect -7 -7 -4 -3
rect -12 -8 -4 -7
rect -12 -12 -11 -8
rect -7 -12 -4 -8
rect -12 -13 -4 -12
rect -12 -17 -11 -13
rect -7 -17 -4 -13
rect -12 -18 -4 -17
rect -12 -22 -11 -18
rect -7 -22 -4 -18
rect -12 -23 -4 -22
rect -12 -27 -11 -23
rect -7 -27 -4 -23
rect -61 -28 -53 -27
rect -61 -32 -60 -28
rect -56 -32 -53 -28
rect -61 -33 -53 -32
rect -61 -37 -60 -33
rect -56 -37 -53 -33
rect -61 -38 -53 -37
rect -61 -42 -60 -38
rect -56 -42 -53 -38
rect -61 -43 -53 -42
rect -61 -47 -60 -43
rect -56 -47 -53 -43
rect -51 -31 -48 -27
rect -44 -31 -43 -27
rect -51 -32 -43 -31
rect -51 -36 -48 -32
rect -44 -36 -43 -32
rect -51 -37 -43 -36
rect -51 -41 -48 -37
rect -44 -41 -43 -37
rect -51 -42 -43 -41
rect -51 -46 -48 -42
rect -44 -46 -43 -42
rect -51 -47 -43 -46
rect -40 -28 -32 -27
rect -40 -32 -39 -28
rect -35 -32 -32 -28
rect -40 -33 -32 -32
rect -40 -37 -39 -33
rect -35 -37 -32 -33
rect -40 -38 -32 -37
rect -40 -42 -39 -38
rect -35 -42 -32 -38
rect -40 -43 -32 -42
rect -40 -47 -39 -43
rect -35 -47 -32 -43
rect -30 -31 -27 -27
rect -23 -31 -22 -27
rect -30 -32 -22 -31
rect -30 -36 -27 -32
rect -23 -36 -22 -32
rect -30 -37 -22 -36
rect -30 -41 -27 -37
rect -23 -41 -22 -37
rect -30 -42 -22 -41
rect -30 -46 -27 -42
rect -23 -46 -22 -42
rect -30 -47 -22 -46
rect -12 -28 -4 -27
rect -12 -32 -11 -28
rect -7 -32 -4 -28
rect -12 -33 -4 -32
rect -12 -37 -11 -33
rect -7 -37 -4 -33
rect -12 -38 -4 -37
rect -12 -42 -11 -38
rect -7 -42 -4 -38
rect -12 -43 -4 -42
rect -12 -47 -11 -43
rect -7 -47 -4 -43
rect -2 9 1 13
rect 5 9 6 13
rect -2 8 6 9
rect -2 4 1 8
rect 5 4 6 8
rect -2 3 6 4
rect -2 -1 1 3
rect 5 -1 6 3
rect -2 -2 6 -1
rect -2 -6 1 -2
rect 5 -6 6 -2
rect -2 -7 6 -6
rect -2 -11 1 -7
rect 5 -11 6 -7
rect -2 -12 6 -11
rect -2 -16 1 -12
rect 5 -16 6 -12
rect -2 -17 6 -16
rect -2 -21 1 -17
rect 5 -21 6 -17
rect -2 -22 6 -21
rect -2 -26 1 -22
rect 5 -26 6 -22
rect -2 -27 6 -26
rect -2 -31 1 -27
rect 5 -31 6 -27
rect -2 -32 6 -31
rect -2 -36 1 -32
rect 5 -36 6 -32
rect -2 -37 6 -36
rect -2 -41 1 -37
rect 5 -41 6 -37
rect -2 -42 6 -41
rect -2 -46 1 -42
rect 5 -46 6 -42
rect -2 -47 6 -46
<< ndcontact >>
rect 3 93 7 97
rect -203 61 -199 65
rect -203 56 -199 60
rect -203 51 -199 55
rect -203 46 -199 50
rect -191 60 -187 64
rect -191 55 -187 59
rect -191 50 -187 54
rect -191 45 -187 49
rect -182 61 -178 65
rect -182 56 -178 60
rect -182 51 -178 55
rect -182 46 -178 50
rect -170 60 -166 64
rect 3 88 7 92
rect 3 83 7 87
rect 3 78 7 82
rect 3 73 7 77
rect 3 68 7 72
rect 3 63 7 67
rect -170 55 -166 59
rect -170 50 -166 54
rect -129 56 -125 60
rect -129 51 -125 55
rect -117 55 -113 59
rect -117 50 -113 54
rect -108 56 -104 60
rect -108 51 -104 55
rect -96 55 -92 59
rect -96 50 -92 54
rect -87 56 -83 60
rect -87 51 -83 55
rect -75 55 -71 59
rect 3 58 7 62
rect -75 50 -71 54
rect -48 53 -44 57
rect -170 45 -166 49
rect -48 48 -44 52
rect -48 43 -44 47
rect -48 38 -44 42
rect -36 52 -32 56
rect -36 47 -32 51
rect -36 42 -32 46
rect -36 37 -32 41
rect -27 51 -23 55
rect -27 46 -23 50
rect -27 41 -23 45
rect -15 52 -11 56
rect -15 47 -11 51
rect -15 42 -11 46
rect -15 37 -11 41
rect 3 53 7 57
rect 3 48 7 52
rect 3 43 7 47
rect 3 38 7 42
rect 15 92 19 96
rect 15 87 19 91
rect 40 95 44 99
rect 40 90 44 94
rect 52 94 56 98
rect 52 89 56 93
rect 61 95 65 99
rect 61 90 65 94
rect 73 94 77 98
rect 73 89 77 93
rect 15 82 19 86
rect 15 77 19 81
rect 15 72 19 76
rect 15 67 19 71
rect 15 62 19 66
rect 15 57 19 61
rect 94 59 98 69
rect 102 59 106 69
rect 110 59 114 69
rect 118 59 122 69
rect 15 52 19 56
rect 15 47 19 51
rect 15 42 19 46
rect 15 37 19 41
rect -187 -6 -183 -2
rect -219 -12 -215 -8
rect -219 -17 -215 -13
rect -219 -22 -215 -18
rect -219 -27 -215 -23
rect -219 -32 -215 -28
rect -219 -37 -215 -33
rect -219 -42 -215 -38
rect -219 -47 -215 -43
rect -219 -52 -215 -48
rect -219 -57 -215 -53
rect -219 -62 -215 -58
rect -219 -67 -215 -63
rect -219 -72 -215 -68
rect -219 -77 -215 -73
rect -219 -82 -215 -78
rect -219 -87 -215 -83
rect -219 -92 -215 -88
rect -219 -97 -215 -93
rect -219 -102 -215 -98
rect -219 -107 -215 -103
rect -207 -13 -203 -9
rect -207 -18 -203 -14
rect -207 -23 -203 -19
rect -187 -11 -183 -7
rect -187 -16 -183 -12
rect -187 -21 -183 -17
rect -175 -7 -171 -3
rect -175 -12 -171 -8
rect -175 -17 -171 -13
rect -175 -22 -171 -18
rect -166 -6 -162 -2
rect -166 -11 -162 -7
rect -166 -16 -162 -12
rect -166 -21 -162 -17
rect -154 -7 -150 -3
rect -154 -12 -150 -8
rect -154 -17 -150 -13
rect -154 -22 -150 -18
rect -207 -28 -203 -24
rect -207 -33 -203 -29
rect -207 -38 -203 -34
rect -207 -43 -203 -39
rect -207 -48 -203 -44
rect 34 1 38 5
rect 34 -4 38 0
rect 46 0 50 4
rect 46 -5 50 -1
rect 55 1 59 5
rect 55 -4 59 0
rect 67 0 71 4
rect 67 -5 71 -1
rect -207 -53 -203 -49
rect -207 -58 -203 -54
rect -207 -63 -203 -59
rect -207 -68 -203 -64
rect -207 -73 -203 -69
rect -207 -78 -203 -74
rect -207 -83 -203 -79
rect -207 -88 -203 -84
rect -60 -73 -56 -69
rect -60 -78 -56 -74
rect -60 -83 -56 -79
rect -60 -88 -56 -84
rect -48 -74 -44 -70
rect -48 -79 -44 -75
rect -48 -84 -44 -80
rect -48 -89 -44 -85
rect -39 -73 -35 -69
rect -39 -78 -35 -74
rect -39 -83 -35 -79
rect -39 -88 -35 -84
rect -27 -74 -23 -70
rect -27 -79 -23 -75
rect -27 -84 -23 -80
rect -27 -89 -23 -85
rect -207 -93 -203 -89
rect -207 -98 -203 -94
rect -207 -103 -203 -99
rect -207 -108 -203 -104
rect -44 -130 -40 -126
rect -44 -135 -40 -131
rect -44 -140 -40 -136
rect -44 -145 -40 -141
rect -32 -131 -28 -127
rect -32 -136 -28 -132
rect -32 -141 -28 -137
rect -32 -146 -28 -142
rect -23 -130 -19 -126
rect -23 -135 -19 -131
rect -23 -140 -19 -136
rect -23 -145 -19 -141
rect -11 -131 -7 -127
rect -11 -136 -7 -132
rect -11 -141 -7 -137
rect -11 -146 -7 -142
<< pdcontact >>
rect -154 142 -150 146
rect -154 137 -150 141
rect -154 132 -150 136
rect -154 127 -150 131
rect -154 122 -150 126
rect -154 117 -150 121
rect -154 112 -150 116
rect -154 107 -150 111
rect -203 102 -199 106
rect -203 97 -199 101
rect -203 92 -199 96
rect -203 87 -199 91
rect -191 103 -187 107
rect -191 98 -187 102
rect -191 93 -187 97
rect -191 88 -187 92
rect -182 102 -178 106
rect -182 97 -178 101
rect -182 92 -178 96
rect -182 87 -178 91
rect -170 103 -166 107
rect -170 98 -166 102
rect -170 93 -166 97
rect -170 88 -166 92
rect -154 102 -150 106
rect -154 97 -150 101
rect -154 92 -150 96
rect -154 87 -150 91
rect -142 143 -138 147
rect -142 138 -138 142
rect 40 139 44 143
rect -142 133 -138 137
rect -142 128 -138 132
rect -142 123 -138 127
rect 40 134 44 138
rect 3 126 7 130
rect -142 118 -138 122
rect -142 113 -138 117
rect -142 108 -138 112
rect -39 117 -35 121
rect -39 112 -35 116
rect -142 103 -138 107
rect -39 107 -35 111
rect -142 98 -138 102
rect -142 93 -138 97
rect -142 88 -138 92
rect -129 100 -125 104
rect -129 95 -125 99
rect -129 90 -125 94
rect -129 85 -125 89
rect -117 101 -113 105
rect -117 96 -113 100
rect -117 91 -113 95
rect -117 86 -113 90
rect -108 100 -104 104
rect -108 95 -104 99
rect -108 90 -104 94
rect -108 85 -104 89
rect -96 101 -92 105
rect -96 96 -92 100
rect -96 91 -92 95
rect -96 86 -92 90
rect -87 100 -83 104
rect -87 95 -83 99
rect -87 90 -83 94
rect -87 85 -83 89
rect -75 101 -71 105
rect -39 102 -35 106
rect -27 118 -23 122
rect -27 113 -23 117
rect 3 121 7 125
rect 3 116 7 120
rect -27 108 -23 112
rect -27 103 -23 107
rect 3 111 7 115
rect 15 127 19 131
rect 15 122 19 126
rect 40 129 44 133
rect 40 124 44 128
rect 52 140 56 144
rect 52 135 56 139
rect 52 130 56 134
rect 52 125 56 129
rect 61 139 65 143
rect 61 134 65 138
rect 61 129 65 133
rect 61 124 65 128
rect 73 140 77 144
rect 73 135 77 139
rect 73 130 77 134
rect 73 125 77 129
rect 15 117 19 121
rect 15 112 19 116
rect -75 96 -71 100
rect -75 91 -71 95
rect -75 86 -71 90
rect 94 107 98 147
rect 107 107 111 147
rect 115 127 119 147
rect -48 84 -44 88
rect -48 79 -44 83
rect -48 74 -44 78
rect -48 69 -44 73
rect -36 85 -32 89
rect -36 80 -32 84
rect -36 75 -32 79
rect -36 70 -32 74
rect -27 84 -23 88
rect -27 79 -23 83
rect -27 74 -23 78
rect -27 69 -23 73
rect -15 85 -11 89
rect -15 80 -11 84
rect -15 75 -11 79
rect -15 70 -11 74
rect 34 45 38 49
rect 34 40 38 44
rect 34 35 38 39
rect 34 30 38 34
rect 46 46 50 50
rect 46 41 50 45
rect 46 36 50 40
rect 46 31 50 35
rect 55 45 59 49
rect 55 40 59 44
rect 55 35 59 39
rect 55 30 59 34
rect 67 46 71 50
rect 67 41 71 45
rect 67 36 71 40
rect 67 31 71 35
rect -11 8 -7 12
rect -11 3 -7 7
rect -11 -2 -7 2
rect -11 -7 -7 -3
rect -11 -12 -7 -8
rect -11 -17 -7 -13
rect -11 -22 -7 -18
rect -11 -27 -7 -23
rect -60 -32 -56 -28
rect -60 -37 -56 -33
rect -60 -42 -56 -38
rect -60 -47 -56 -43
rect -48 -31 -44 -27
rect -48 -36 -44 -32
rect -48 -41 -44 -37
rect -48 -46 -44 -42
rect -39 -32 -35 -28
rect -39 -37 -35 -33
rect -39 -42 -35 -38
rect -39 -47 -35 -43
rect -27 -31 -23 -27
rect -27 -36 -23 -32
rect -27 -41 -23 -37
rect -27 -46 -23 -42
rect -11 -32 -7 -28
rect -11 -37 -7 -33
rect -11 -42 -7 -38
rect -11 -47 -7 -43
rect 1 9 5 13
rect 1 4 5 8
rect 1 -1 5 3
rect 1 -6 5 -2
rect 1 -11 5 -7
rect 1 -16 5 -12
rect 1 -21 5 -17
rect 1 -26 5 -22
rect 1 -31 5 -27
rect 1 -36 5 -32
rect 1 -41 5 -37
rect 1 -46 5 -42
<< psubstratepcontact >>
rect 34 79 38 83
rect 42 79 46 83
rect 50 79 54 83
rect 59 79 63 83
rect 67 79 71 83
rect 75 79 79 83
rect -56 27 -52 31
rect -48 27 -44 31
rect -40 27 -36 31
rect -32 27 -28 31
rect -24 27 -20 31
rect -16 27 -12 31
rect -8 27 -4 31
rect 0 27 4 31
rect -226 -160 -222 -156
rect -218 -160 -214 -156
rect -210 -160 -206 -156
rect -202 -160 -198 -156
rect -194 -160 -190 -156
rect -186 -160 -182 -156
rect -178 -160 -174 -156
rect -170 -160 -166 -156
rect -162 -160 -158 -156
rect -154 -160 -150 -156
rect -146 -160 -142 -156
rect -135 -160 -131 -156
rect -127 -160 -123 -156
rect -119 -160 -115 -156
rect -110 -160 -106 -156
rect -102 -160 -98 -156
rect -93 -160 -89 -156
rect -85 -160 -81 -156
rect -43 -160 -39 -156
rect -35 -160 -31 -156
rect -27 -160 -23 -156
rect -19 -160 -15 -156
rect -11 -160 -7 -156
rect -3 -160 1 -156
rect 28 -160 32 -156
rect 36 -160 40 -156
rect 44 -160 48 -156
rect 53 -160 57 -156
rect 61 -160 65 -156
rect 69 -160 73 -156
rect 90 -159 94 -155
rect 106 -159 110 -155
<< nsubstratencontact >>
rect -203 151 -199 155
rect -195 151 -191 155
rect -187 151 -183 155
rect -179 151 -175 155
rect -171 151 -167 155
rect -163 151 -159 155
rect -155 151 -151 155
rect -147 151 -143 155
rect -139 151 -135 155
rect -126 151 -122 155
rect -118 151 -114 155
rect -109 151 -105 155
rect -101 151 -97 155
rect -93 151 -89 155
rect -84 151 -80 155
rect -76 151 -72 155
rect 35 151 39 155
rect 43 151 47 155
rect 51 151 55 155
rect 60 151 64 155
rect 68 151 72 155
rect 76 151 80 155
rect 90 151 94 155
rect 106 151 110 155
rect -328 141 -316 147
rect -328 5 -316 11
rect -306 141 -294 147
rect -306 5 -294 11
rect -284 139 -272 145
rect -284 3 -272 9
rect -262 141 -250 147
rect -262 5 -250 11
rect -240 141 -228 147
rect -240 5 -228 11
rect -45 139 -41 143
rect -37 139 -33 143
rect -29 139 -25 143
rect -21 139 -17 143
rect -13 139 -9 143
rect -5 139 -1 143
rect 3 139 7 143
rect 11 139 15 143
rect 29 56 33 60
rect 37 56 41 60
rect 45 56 49 60
rect 54 56 58 60
rect 62 56 66 60
rect -60 17 -56 21
rect -52 17 -48 21
rect -44 17 -40 21
rect -36 17 -32 21
rect -28 17 -24 21
rect -20 17 -16 21
rect -12 17 -8 21
rect -4 17 0 21
rect 4 17 8 21
<< polysilicon >>
rect -147 147 -145 150
rect 99 147 101 149
rect 104 147 106 149
rect 112 147 114 149
rect -196 107 -194 110
rect -175 107 -173 110
rect 47 144 49 147
rect 68 144 70 147
rect -32 134 12 136
rect -32 122 -30 134
rect 10 131 12 134
rect -122 105 -120 108
rect -101 105 -99 108
rect -80 105 -78 108
rect -196 82 -194 87
rect -175 82 -173 87
rect -147 79 -145 87
rect 10 108 12 111
rect -32 101 -30 102
rect -52 97 -30 101
rect -41 89 -39 92
rect -20 89 -18 108
rect 10 97 12 100
rect 47 99 49 124
rect 68 99 70 124
rect 112 126 114 127
rect 112 124 117 126
rect -196 65 -194 68
rect -175 65 -173 70
rect -122 60 -120 85
rect -101 60 -99 85
rect -80 60 -78 85
rect -41 67 -39 69
rect -51 65 -39 67
rect -20 66 -18 69
rect -41 57 -39 58
rect -20 57 -18 58
rect -122 47 -120 50
rect -101 47 -99 50
rect -80 47 -78 50
rect -196 40 -194 45
rect -175 42 -173 45
rect 47 86 49 89
rect 68 86 70 89
rect 99 76 101 107
rect 104 96 106 107
rect 104 94 109 96
rect 107 86 109 94
rect 98 72 101 76
rect 99 69 101 72
rect 107 69 109 82
rect 115 69 117 124
rect 99 57 101 59
rect 107 57 109 59
rect 115 57 117 59
rect 41 50 43 53
rect 62 50 64 53
rect -41 34 -39 37
rect -20 34 -18 37
rect 10 34 12 37
rect -4 13 -2 16
rect -180 -2 -178 9
rect -159 -2 -157 9
rect -212 -8 -210 -5
rect -180 -25 -178 -22
rect -159 -25 -157 -22
rect -53 -27 -51 -24
rect -32 -27 -30 -24
rect 41 5 43 30
rect 62 5 64 30
rect 41 -8 43 -5
rect 62 -8 64 -5
rect -53 -52 -51 -47
rect -32 -52 -30 -47
rect -4 -55 -2 -47
rect -53 -69 -51 -66
rect -32 -69 -30 -64
rect -53 -94 -51 -89
rect -32 -92 -30 -89
rect -212 -111 -210 -108
rect -37 -126 -35 -115
rect -16 -126 -14 -115
rect -37 -149 -35 -146
rect -16 -149 -14 -146
<< polycontact >>
rect -196 78 -192 82
rect -177 78 -173 82
rect -20 108 -16 112
rect -56 97 -52 101
rect 8 100 12 104
rect 43 103 47 107
rect 64 103 68 107
rect -145 79 -141 83
rect -177 70 -173 74
rect -126 64 -122 68
rect -105 64 -101 68
rect -84 64 -80 68
rect -55 63 -51 67
rect -41 58 -37 62
rect -22 58 -18 62
rect -80 43 -76 47
rect -196 36 -192 40
rect 111 100 115 104
rect 106 82 110 86
rect 94 72 98 76
rect -180 9 -176 13
rect -161 9 -157 13
rect -212 -5 -208 -1
rect -159 -29 -155 -25
rect 37 9 41 13
rect 58 9 62 13
rect -53 -56 -49 -52
rect -34 -56 -30 -52
rect -2 -55 2 -51
rect -34 -64 -30 -60
rect -53 -98 -49 -94
rect -37 -115 -33 -111
rect -18 -115 -14 -111
<< metal1 >>
rect -220 156 -216 158
rect -328 152 -309 156
rect -328 147 -316 152
rect -328 -4 -316 5
rect -313 0 -309 152
rect -306 152 -287 156
rect -306 147 -294 152
rect -306 0 -294 5
rect -313 -4 -294 0
rect -291 0 -287 152
rect -284 150 -265 154
rect -284 145 -272 150
rect -284 0 -272 3
rect -291 -4 -272 0
rect -269 0 -265 150
rect -262 152 -243 156
rect -262 147 -250 152
rect -262 0 -250 5
rect -269 -4 -250 0
rect -247 0 -243 152
rect -240 155 126 156
rect -240 151 -203 155
rect -199 151 -195 155
rect -191 151 -187 155
rect -183 151 -179 155
rect -175 151 -171 155
rect -167 151 -163 155
rect -159 151 -155 155
rect -151 151 -147 155
rect -143 151 -139 155
rect -135 151 -126 155
rect -122 151 -118 155
rect -114 151 -109 155
rect -105 151 -101 155
rect -97 151 -93 155
rect -89 151 -84 155
rect -80 151 -76 155
rect -72 151 35 155
rect 39 151 43 155
rect 47 151 51 155
rect 55 151 60 155
rect 64 151 68 155
rect 72 151 76 155
rect 80 151 90 155
rect 94 151 106 155
rect 110 151 126 155
rect -240 150 126 151
rect -240 147 -228 150
rect -203 106 -199 150
rect -240 0 -228 5
rect -220 0 -216 101
rect -203 101 -199 102
rect -203 96 -199 97
rect -203 91 -199 92
rect -191 102 -187 103
rect -191 97 -187 98
rect -191 92 -187 93
rect -191 82 -187 88
rect -182 106 -178 150
rect -154 146 -150 150
rect -154 141 -150 142
rect -154 136 -150 137
rect -154 131 -150 132
rect -154 126 -150 127
rect -154 121 -150 122
rect -154 116 -150 117
rect -154 111 -150 112
rect -182 101 -178 102
rect -182 96 -178 97
rect -182 91 -178 92
rect -170 102 -166 103
rect -170 97 -166 98
rect -170 92 -166 93
rect -192 78 -177 82
rect -203 60 -199 61
rect -203 55 -199 56
rect -203 50 -199 51
rect -211 46 -203 49
rect -211 45 -199 46
rect -191 64 -187 78
rect -170 77 -166 88
rect -154 106 -150 107
rect -154 101 -150 102
rect -154 96 -150 97
rect -154 91 -150 92
rect -142 142 -138 143
rect -142 137 -138 138
rect -142 132 -138 133
rect -142 127 -138 128
rect -142 122 -138 123
rect -142 117 -138 118
rect -142 112 -138 113
rect -142 107 -138 108
rect -142 102 -138 103
rect -142 97 -138 98
rect -142 92 -138 93
rect -129 104 -125 150
rect -129 99 -125 100
rect -129 94 -125 95
rect -138 88 -133 92
rect -184 70 -181 74
rect -145 77 -141 79
rect -191 59 -187 60
rect -191 54 -187 55
rect -191 49 -187 50
rect -182 60 -178 61
rect -182 55 -178 56
rect -182 50 -178 51
rect -211 30 -207 45
rect -182 30 -178 46
rect -170 64 -166 73
rect -137 68 -133 88
rect -129 89 -125 90
rect -117 100 -113 101
rect -117 95 -113 96
rect -117 90 -113 91
rect -117 68 -113 86
rect -108 104 -104 150
rect -108 99 -104 100
rect -108 94 -104 95
rect -108 89 -104 90
rect -96 100 -92 101
rect -96 95 -92 96
rect -96 90 -92 91
rect -96 68 -92 86
rect -87 104 -83 150
rect -64 139 -45 143
rect -41 139 -37 143
rect -33 139 -29 143
rect -25 139 -21 143
rect -17 139 -13 143
rect -9 139 -5 143
rect -1 139 3 143
rect 7 139 11 143
rect 15 139 19 143
rect -87 99 -83 100
rect -87 94 -83 95
rect -87 89 -83 90
rect -75 100 -71 101
rect -75 95 -71 96
rect -75 90 -71 91
rect -75 68 -71 86
rect -64 68 -60 139
rect -39 121 -35 139
rect 3 130 7 139
rect 3 125 7 126
rect -39 116 -35 117
rect -39 111 -35 112
rect -39 106 -35 107
rect -27 117 -23 118
rect -27 112 -23 113
rect 3 120 7 121
rect 3 115 7 116
rect 15 126 19 127
rect 15 121 19 122
rect 15 116 19 117
rect -27 107 -23 108
rect 15 107 19 112
rect -27 96 -23 103
rect -48 92 -23 96
rect -48 88 -44 92
rect -48 83 -44 84
rect -48 78 -44 79
rect -48 73 -44 74
rect -36 84 -32 85
rect -36 79 -32 80
rect -36 74 -32 75
rect -170 59 -166 60
rect -170 54 -166 55
rect -170 49 -166 50
rect -154 64 -126 68
rect -117 64 -105 68
rect -96 64 -84 68
rect -75 64 -60 68
rect -211 26 -175 30
rect -247 -4 -228 0
rect -221 -1 -216 0
rect -207 9 -192 13
rect -188 9 -180 13
rect -176 9 -161 13
rect -207 -1 -203 9
rect -221 -4 -212 -1
rect -220 -5 -212 -4
rect -208 -5 -203 -1
rect -219 -13 -215 -12
rect -219 -18 -215 -17
rect -219 -23 -215 -22
rect -219 -28 -215 -27
rect -219 -33 -215 -32
rect -219 -38 -215 -37
rect -219 -43 -215 -42
rect -219 -48 -215 -47
rect -219 -53 -215 -52
rect -219 -58 -215 -57
rect -219 -63 -215 -62
rect -219 -68 -215 -67
rect -219 -73 -215 -72
rect -219 -78 -215 -77
rect -219 -83 -215 -82
rect -219 -88 -215 -87
rect -219 -93 -215 -92
rect -219 -98 -215 -97
rect -219 -103 -215 -102
rect -219 -154 -215 -107
rect -207 -9 -203 -5
rect -207 -14 -203 -13
rect -207 -19 -203 -18
rect -207 -24 -203 -23
rect -207 -29 -203 -28
rect -207 -34 -203 -33
rect -207 -39 -203 -38
rect -207 -44 -203 -43
rect -207 -49 -203 -48
rect -207 -54 -203 -53
rect -207 -59 -203 -58
rect -207 -64 -203 -63
rect -207 -69 -203 -68
rect -207 -74 -203 -73
rect -207 -79 -203 -78
rect -207 -84 -203 -83
rect -207 -89 -203 -88
rect -207 -94 -203 -93
rect -207 -99 -203 -98
rect -207 -104 -203 -103
rect -187 -7 -183 -6
rect -187 -12 -183 -11
rect -187 -17 -183 -16
rect -187 -154 -183 -21
rect -175 -3 -171 -1
rect -175 -8 -171 -7
rect -175 -13 -171 -12
rect -175 -18 -171 -17
rect -166 -7 -162 -6
rect -166 -12 -162 -11
rect -166 -17 -162 -16
rect -166 -154 -162 -21
rect -154 -3 -150 64
rect -154 -8 -150 -7
rect -154 -13 -150 -12
rect -154 -18 -150 -17
rect -129 55 -125 56
rect -155 -111 -151 -25
rect -129 -154 -125 51
rect -117 59 -113 64
rect -117 54 -113 55
rect -108 55 -104 56
rect -108 -154 -104 51
rect -96 59 -92 64
rect -96 54 -92 55
rect -87 55 -83 56
rect -87 31 -83 51
rect -75 59 -71 64
rect -75 54 -71 55
rect -87 -154 -83 27
rect -76 21 -72 47
rect -55 41 -51 63
rect -36 62 -32 70
rect -27 88 -23 92
rect -27 83 -23 84
rect -27 78 -23 79
rect -27 73 -23 74
rect -15 100 8 104
rect -15 89 -11 100
rect -15 84 -11 85
rect -15 79 -11 80
rect -15 74 -11 75
rect -37 58 -22 62
rect -48 52 -44 53
rect -48 47 -44 48
rect -48 42 -44 43
rect -48 31 -44 38
rect -36 56 -32 58
rect -15 56 -11 70
rect -36 51 -32 52
rect -36 46 -32 47
rect -36 41 -32 42
rect -27 50 -23 51
rect -27 45 -23 46
rect -27 31 -23 41
rect -15 51 -11 52
rect -15 46 -11 47
rect -15 41 -11 42
rect 3 92 7 93
rect 3 87 7 88
rect 3 82 7 83
rect 3 77 7 78
rect 3 72 7 73
rect 3 67 7 68
rect 3 62 7 63
rect 3 57 7 58
rect 3 52 7 53
rect 3 47 7 48
rect 3 42 7 43
rect 3 31 7 38
rect 15 96 19 103
rect 15 91 19 92
rect 15 86 19 87
rect 15 81 19 82
rect 15 76 19 77
rect 15 71 19 72
rect 15 66 19 67
rect 15 61 19 62
rect 15 56 19 57
rect 24 60 28 150
rect 40 143 44 150
rect 40 138 44 139
rect 40 133 44 134
rect 40 128 44 129
rect 52 139 56 140
rect 52 134 56 135
rect 52 129 56 130
rect 52 107 56 125
rect 61 143 65 150
rect 107 147 111 150
rect 61 138 65 139
rect 61 133 65 134
rect 61 128 65 129
rect 73 139 77 140
rect 73 134 77 135
rect 73 129 77 130
rect 41 103 43 107
rect 52 103 64 107
rect 40 94 44 95
rect 40 83 44 90
rect 52 98 56 103
rect 52 93 56 94
rect 61 94 65 95
rect 61 83 65 90
rect 73 98 77 125
rect 116 124 122 127
rect 94 104 98 107
rect 94 101 111 104
rect 73 93 77 94
rect 77 89 106 93
rect 111 92 114 100
rect 119 97 122 124
rect 119 93 124 97
rect 111 89 116 92
rect 33 79 34 83
rect 38 79 42 83
rect 46 79 50 83
rect 54 79 59 83
rect 63 79 67 83
rect 71 79 75 83
rect 79 79 83 83
rect 102 82 106 89
rect 113 77 116 89
rect 72 72 94 76
rect 103 74 116 77
rect 24 56 29 60
rect 33 56 37 60
rect 41 56 45 60
rect 49 56 54 60
rect 58 56 62 60
rect 66 56 68 60
rect 15 51 19 52
rect 15 46 19 47
rect 15 41 19 42
rect 34 49 38 56
rect 34 44 38 45
rect 34 39 38 40
rect 34 34 38 35
rect -59 27 -56 31
rect -52 27 -48 31
rect -44 27 -40 31
rect -36 27 -32 31
rect -28 27 -24 31
rect -20 27 -16 31
rect -12 27 -8 31
rect -4 27 0 31
rect 4 27 10 31
rect 46 45 50 46
rect 46 40 50 41
rect 46 35 50 36
rect -76 17 -60 21
rect -56 17 -52 21
rect -48 17 -44 21
rect -40 17 -36 21
rect -32 17 -28 21
rect -24 17 -20 21
rect -16 17 -12 21
rect -8 17 -4 21
rect 0 17 4 21
rect 8 17 10 21
rect -60 -28 -56 17
rect -60 -33 -56 -32
rect -60 -38 -56 -37
rect -60 -43 -56 -42
rect -48 -32 -44 -31
rect -48 -37 -44 -36
rect -48 -42 -44 -41
rect -48 -52 -44 -46
rect -39 -28 -35 17
rect -11 12 -7 17
rect 46 13 50 31
rect 55 49 59 56
rect 72 50 76 72
rect 103 69 106 74
rect 119 69 122 93
rect 94 56 98 59
rect 87 52 98 56
rect 55 44 59 45
rect 55 39 59 40
rect 55 34 59 35
rect 71 46 76 50
rect 67 45 71 46
rect 67 40 71 41
rect 67 35 71 36
rect -11 7 -7 8
rect -11 2 -7 3
rect -11 -3 -7 -2
rect -11 -8 -7 -7
rect -11 -13 -7 -12
rect -11 -18 -7 -17
rect -11 -23 -7 -22
rect -39 -33 -35 -32
rect -39 -38 -35 -37
rect -39 -43 -35 -42
rect -27 -32 -23 -31
rect -27 -37 -23 -36
rect -27 -42 -23 -41
rect -49 -56 -34 -52
rect -60 -74 -56 -73
rect -60 -79 -56 -78
rect -60 -84 -56 -83
rect -68 -88 -60 -85
rect -68 -89 -56 -88
rect -48 -70 -44 -56
rect -27 -57 -23 -46
rect -11 -28 -7 -27
rect -11 -33 -7 -32
rect -11 -38 -7 -37
rect -11 -43 -7 -42
rect 5 9 37 13
rect 46 9 58 13
rect 1 8 5 9
rect 1 3 5 4
rect 1 -2 5 -1
rect 1 -7 5 -6
rect 1 -12 5 -11
rect 1 -17 5 -16
rect 1 -22 5 -21
rect 1 -27 5 -26
rect 1 -32 5 -31
rect 1 -37 5 -36
rect 1 -42 5 -41
rect 34 0 38 1
rect 5 -46 10 -42
rect -2 -57 2 -55
rect -48 -75 -44 -74
rect -48 -80 -44 -79
rect -48 -85 -44 -84
rect -39 -74 -35 -73
rect -39 -79 -35 -78
rect -39 -84 -35 -83
rect -68 -104 -64 -89
rect -45 -98 -42 -94
rect -39 -104 -35 -88
rect -27 -70 -23 -61
rect 6 -66 10 -46
rect -27 -75 -23 -74
rect -27 -80 -23 -79
rect -27 -85 -23 -84
rect -11 -70 10 -66
rect -68 -108 -32 -104
rect -66 -115 -37 -111
rect -33 -115 -18 -111
rect -44 -131 -40 -130
rect -44 -136 -40 -135
rect -44 -141 -40 -140
rect -44 -154 -40 -145
rect -32 -127 -28 -125
rect -32 -132 -28 -131
rect -32 -137 -28 -136
rect -32 -142 -28 -141
rect -23 -131 -19 -130
rect -23 -136 -19 -135
rect -23 -141 -19 -140
rect -23 -154 -19 -145
rect -11 -127 -7 -70
rect -11 -132 -7 -131
rect -11 -137 -7 -136
rect -11 -142 -7 -141
rect 34 -154 38 -4
rect 46 4 50 9
rect 46 -1 50 0
rect 55 0 59 1
rect 55 -154 59 -4
rect 67 4 71 31
rect 67 -1 71 0
rect 94 -154 98 52
rect 110 -154 114 59
rect -229 -155 126 -154
rect -229 -156 90 -155
rect -229 -160 -226 -156
rect -222 -160 -218 -156
rect -214 -160 -210 -156
rect -206 -160 -202 -156
rect -198 -160 -194 -156
rect -190 -160 -186 -156
rect -182 -160 -178 -156
rect -174 -160 -170 -156
rect -166 -160 -162 -156
rect -158 -160 -154 -156
rect -150 -160 -146 -156
rect -142 -160 -135 -156
rect -131 -160 -127 -156
rect -123 -160 -119 -156
rect -115 -160 -110 -156
rect -106 -160 -102 -156
rect -98 -160 -93 -156
rect -89 -160 -85 -156
rect -81 -160 -43 -156
rect -39 -160 -35 -156
rect -31 -160 -27 -156
rect -23 -160 -19 -156
rect -15 -160 -11 -156
rect -7 -160 -3 -156
rect 1 -160 28 -156
rect 32 -160 36 -156
rect 40 -160 44 -156
rect 48 -160 53 -156
rect 57 -160 61 -156
rect 65 -160 69 -156
rect 73 -159 90 -156
rect 94 -159 106 -155
rect 110 -159 126 -155
rect 73 -160 126 -159
<< m2contact >>
rect -332 -4 -328 0
rect -220 101 -216 105
rect -181 70 -177 74
rect -170 73 -166 77
rect -145 73 -141 77
rect -192 36 -188 40
rect -56 101 -52 105
rect -16 108 -12 112
rect -175 26 -171 30
rect -225 -4 -221 0
rect -192 9 -188 13
rect -175 -1 -171 3
rect -155 -115 -151 -111
rect -87 27 -83 31
rect 15 103 19 107
rect -55 37 -51 41
rect 37 103 41 107
rect 83 79 87 83
rect -63 27 -59 31
rect 83 52 87 56
rect -38 -64 -34 -60
rect -27 -61 -23 -57
rect -2 -61 2 -57
rect -49 -98 -45 -94
rect -32 -108 -28 -104
rect -70 -115 -66 -111
rect -32 -125 -28 -121
<< metal2 >>
rect -48 108 -16 112
rect -216 101 -56 105
rect -166 73 -145 77
rect -181 64 -177 70
rect -48 64 -44 108
rect -181 60 -44 64
rect -192 13 -188 36
rect -83 27 -63 31
rect -175 3 -171 26
rect -328 -4 -225 0
rect -55 -59 -51 37
rect -55 -63 -45 -59
rect -49 -94 -45 -63
rect -38 -60 -34 108
rect 19 103 37 107
rect 83 56 87 79
rect -23 -61 -2 -57
rect -151 -115 -70 -111
rect -32 -121 -28 -108
<< pseudo_rnwell >>
rect -329 147 -315 148
rect -329 5 -328 147
rect -316 5 -315 147
rect -329 4 -315 5
rect -307 147 -293 148
rect -307 5 -306 147
rect -294 5 -293 147
rect -263 147 -249 148
rect -307 4 -293 5
rect -285 145 -271 146
rect -285 3 -284 145
rect -272 3 -271 145
rect -263 5 -262 147
rect -250 5 -249 147
rect -263 4 -249 5
rect -241 147 -227 148
rect -241 5 -240 147
rect -228 5 -227 147
rect -241 4 -227 5
rect -285 2 -271 3
<< rnwell >>
rect -328 11 -316 141
rect -306 11 -294 141
rect -284 9 -272 139
rect -262 11 -250 141
rect -240 11 -228 141
<< labels >>
rlabel metal1 123 95 123 95 1 OUT
rlabel metal1 -228 -158 -228 -158 1 0
rlabel metal1 -183 72 -183 72 1 INP
rlabel metal1 -44 -96 -44 -96 1 INN
rlabel metal1 -218 157 -218 157 5 En
<< end >>
